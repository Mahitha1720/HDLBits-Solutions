//Description: The output is assigned the value to be same as the input

module top_module( input in, output out );
   assign out=in;
endmodule
