//Description: The AND gate-level logic is implemented

module top_module( 
    input a, 
    input b, 
    output out );
    assign out=a&b;
endmodule
