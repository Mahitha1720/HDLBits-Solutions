// Description: Output constant logic 1

module top_module(
    output one
);

  // Output is given to be high i.e. 1
assign one = 1'b1;

endmodule
