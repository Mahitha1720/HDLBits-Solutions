module top_module( 
    input [399:0] a, b,
    input cin,
    output cout,
    output [399:0] sum
);

    genvar i;
    wire[99:0] w;
	
    generate
        bcd_fadd(a[3:0], b[3:0], cin, w[0],sum[3:0]);
        for (i=4; i<400; i=i+4)
			begin: bcd_adder
				bcd_fadd bcd_adder(a[i+3:i], b[i+3:i], w[i/4-1],w[i/4],sum[i+3:i]);
			end
    endgenerate
    
    assign cout = w[99];
	
endmodule
