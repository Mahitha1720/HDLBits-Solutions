//Description: Creating a NOT gate, where output is complement of input

module top_module( input in, output out );
   assign out=~in;
endmodule
