//Description:No input and output is hardwired to be zero


module top_module(
    output zero
);

    assign zero = 1'b0;

endmodule
